`timescale 1ns / 1ps

module instr_mem(PC, Instr);

    input [31:0] PC;
    output wire [31:0] Instr;

    reg [31:0] RAM[63:0];

    initial begin  // Copy of instructions found on page 453.
        RAM[ 0] <= 32'b11100000010011110000000000001111;
        RAM[ 1] <= 32'b11100010100000000010000000000101;
        RAM[ 2] <= 32'b11100010100000000011000000001100;
        RAM[ 3] <= 32'b11100010010000110111000000001001;
        RAM[ 4] <= 32'b11100001100001110100000000000010;
        RAM[ 5] <= 32'b11100000000000110101000000000100;
        RAM[ 6] <= 32'b11100000100001010101000000000100;
        RAM[ 7] <= 32'b11100000010101011000000000000111;
        RAM[ 8] <= 32'b00001010000000000000000000001100;
        RAM[ 9] <= 32'b11100000010100111000000000000100;
        RAM[10] <= 32'b10101010000000000000000000000000;
        RAM[11] <= 32'b11100010100000000101000000000000;
        RAM[12] <= 32'b11100000010101111000000000000010;
        RAM[13] <= 32'b10110010100001010111000000000001;
        RAM[14] <= 32'b11100000010001110111000000000010;
        RAM[15] <= 32'b11100101100000110111000001010100;
        RAM[16] <= 32'b11100101100100000010000001100000;
        RAM[17] <= 32'b11100000100011111111000000000000;
        RAM[18] <= 32'b11100010100000000010000000000001;
        RAM[19] <= 32'b11101010000000000000000000000001;
        RAM[20] <= 32'b11100010100000000010000000000001;
        RAM[21] <= 32'b11100010100000000010000000000001;
        RAM[22] <= 32'b11100101100000000010000001010100;
    end

    assign Instr = RAM[PC[31:2]];  // 2 here because we want to word align mem read.

endmodule

