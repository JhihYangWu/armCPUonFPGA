`timescale 1ns / 1ps

module mux8x1_tb();

    reg [31:0] A0, A1, A2, A3, A4, A5, A6, A7;
    reg [2:0] select;
    wire [31:0] Y;

    mux8x1 a1(A0, A1, A2, A3, A4, A5, A6, A7, select, Y);

    initial begin
        select <= 0; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 1; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 2; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 3; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 4; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 5; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 6; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 7; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 6; #100;
        select <= 7; A0 <= 12; A1 <= 31; A2 <= 45; A3 <= 121; A4 <= 1234; A5 <= 21312; A6 <= 1; A7 <= 3123; #100;

    end

endmodule

