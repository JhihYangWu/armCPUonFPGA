`timescale 1ns / 1ps

module comparator_tb();

    reg [31:0] A, B;
    wire eq, neq, lt, lte, gt, gte;

    comparator #(32) a1(A, B, eq, neq, lt, lte, gt, gte);

    initial begin
        A <= 0; B <= 0; #100;
        A <= 2648; B <= 5357; #100;
        A <= 967; B <= 4448; #100;
        A <= 3207; B <= 7360; #100;
        A <= 787; B <= 1735; #100;
        A <= 4300; B <= 7550; #100;
        A <= 9874; B <= 9875; #100;
        A <= 5580; B <= 5579; #100;
        A <= 9425; B <= 8571; #100;
        A <= 7433; B <= 7433; #100;
        A <= 9488; B <= 4985; #100;
        A <= 7636; B <= 9064; #100;
        A <= 8824; B <= 9435; #100;
        A <= 8344; B <= 7538; #100;
        A <= 4019; B <= 5959; #100;
        A <= 4179; B <= 9270; #100;
        A <= 6636; B <= 1260; #100;
        A <= 2291; B <= 3950; #100;
        A <= 3589; B <= 5637; #100;
        A <= 8714; B <= 8662; #100;
        A <= 3212; B <= 537; #100;
        A <= 6282; B <= 6047; #100;
        A <= 5946; B <= 187; #100;
        A <= 6576; B <= 1136; #100;
        A <= 4843; B <= 2520; #100;
        A <= 1609; B <= 1737; #100;
        A <= 8450; B <= 9990; #100;
        A <= 5521; B <= 2105; #100;

    end

endmodule

